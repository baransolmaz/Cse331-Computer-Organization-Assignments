module and32(in1,in2,result);
	input [31:0] in1,in2;
	output [31:0] result;
	
	and(result[0],in1[0],in2[0]);
	and(result[1],in1[1],in2[1]);
	and(result[2],in1[2],in2[2]);
	and(result[3],in1[3],in2[3]);
	and(result[4],in1[4],in2[4]);
	and(result[5],in1[5],in2[5]);
	and(result[6],in1[6],in2[6]);
	and(result[7],in1[7],in2[7]);
	and(result[8],in1[8],in2[8]);
	and(result[9],in1[9],in2[9]);
	and(result[10],in1[10],in2[10]);
	and(result[11],in1[11],in2[11]);
	and(result[12],in1[12],in2[12]);
	and(result[13],in1[13],in2[13]);
	and(result[14],in1[14],in2[14]);
	and(result[15],in1[15],in2[15]);
	and(result[16],in1[16],in2[16]);
	and(result[17],in1[17],in2[17]);
	and(result[18],in1[18],in2[18]);
	and(result[19],in1[19],in2[19]);
	and(result[20],in1[20],in2[20]);
	and(result[21],in1[21],in2[21]);
	and(result[22],in1[22],in2[22]);
	and(result[23],in1[23],in2[23]);
	and(result[24],in1[24],in2[24]);
	and(result[25],in1[25],in2[25]);
	and(result[26],in1[26],in2[26]);
	and(result[27],in1[27],in2[27]);
	and(result[28],in1[28],in2[28]);
	and(result[29],in1[29],in2[29]);
	and(result[30],in1[30],in2[30]);
	and(result[31],in1[31],in2[31]);
	
endmodule